`ifdef simulation 
    parameter DIV1 = 3;
`else
    parameter DIV1 = 10;
`endif
parameter DIV2 = 5;
