
module issp (
	probe,
	source,
	source_clk);	

	input	[0:0]	probe;
	output	[2:0]	source;
	input		source_clk;
endmodule
