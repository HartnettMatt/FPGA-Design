module aud (
  input wire clk
  );

endmodule // aud
