module aud (
  input clk,
  input reset_n,
  input adcdat,
  inout adclrck,
  inout bclk,
  output dacdat,
  inout daclrck,
  output xck
  );

endmodule // aud
