parameter 
