parameter Wait_STATE    =     4'b0000;
parameter Start_STATE   =     4'b0001;
parameter Address_STATE =     4'b0010;
parameter Ack1_STATE    =     4'b0011;
parameter Data1_STATE   =     4'b0100;
parameter Ack2_STATE    =     4'b0101;
parameter Data2_STATE   =     4'b0110;
parameter Ack3_STATE    =     4'b0111;
parameter Stop_STATE    =     4'b1000;
