`ifdef lowRes
  parameter fPorchH = 16;
  parameter bPorchH = 48;
  parameter dispTimeH = 640;
  parameter pulseWidthH = 96;
  parameter syncTimeH = 800;
`else

`endif
