
module issp1 (
	probe,
	source);	

	input	[5:0]	probe;
	output	[1:0]	source;
endmodule
