module VTC(
  input wire       clock_in,
  output           vSync,
  output           hSync,
  output           hPixel,
  output           line,
  output           video_active
);

endmodule
