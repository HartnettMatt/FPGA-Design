`ifdef lowRes
  parameter fPorchH = 16;
  parameter bPorchH = 48;
  parameter dispTimeH = 640;
  parameter pulseWidthH = 96;
  parameter syncTimeH = 800;
  parameter fPorchV = 10;
  parameter bPorchV = 29;
  parameter dispTimeV = 480;
  parameter pulseWidthV = 2;
  parameter syncTimeV = 521;
`else

`endif
