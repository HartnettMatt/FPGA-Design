module i2c_OL ();
`include "i2c_states.vh"
endmodule // i2c_OL
